module aaa();
	input clk,
	output clk_20
endmodule
